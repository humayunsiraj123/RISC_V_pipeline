module risc_v_pipeline();





endmodule : risc_v_pipeline