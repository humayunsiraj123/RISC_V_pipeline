module register();
endmodule
